Circuito_t2_2

R1 1 2 1.049124789255k
R2 3 2 2.057037410185k
R3 2 5 3.145866332601k
R4 5 1 4.120366732090k
R5 5 6 3.092796241346k
R6 1 4 2.078623037946k
R7 7 8 1.047211798510k


*Independent Sources

Vx 6 8 DC 8.7098

V3 4 7 DC 0

*Dependent Sources

Gb 6 3 2 5 7.2690889775598m
Hc 5 8 V3 8.04305881912k

.control
 op
 print all
 .endc
 .end
