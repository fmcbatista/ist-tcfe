Circuito_t2.2

.INCLUDE ngspice_2.txt

.control
 op
 print all
 .endc
 .end
