Circuito Teste

.options savecurrents

 Va 0 3 5.13416
 R1 1 0 1.0491248k
 R2 2 1 2.0570374k
 R3 1 4 3.1458663k
 R4 3 4 4.1203667k
 R5 4 5 3.0927962k
 R6 3 6 2.0786230k
 R7 aux 7 1.0472118k
 I  7 5 1.0310985m
 Gi 5 2 (1,4) 7.2690898m
 Vctl 6 aux 0
 H1 4 7 Vctl 8.0430588k
 
 .control
 
 op
 
 echo "****************"
 echo "Operating Point"
 echo "****************"
 
 
 echo "op_TAB"
 echo "@Id[i]=1.0311e-3"
 print all
 echo "op_END"
 quit
 .endc
 .end
