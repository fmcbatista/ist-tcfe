Circuit_t2.4

.options savecurrents

.INCLUDE ngspice_4.txt


.ic v(6)=8.7098  v(8)=0

.end

.control



op

echo "Transient Analysis"

tran 1e-6 20ms

plot v(6) v(1)

hardcopy trans.ps v(6) v(1)


.endc


.end
