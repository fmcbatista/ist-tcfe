Circuito_t2

.INCLUDE ngspice_values.txt






.control
 op
 
 echo "Operating Point Analysis"
 
 print  V(6)-V(8) > Vx_p2.txt
 echo "Ia"
 print (v(2)-v(1))/1.0491248k
 echo "ib"
 print (v(3)-v(2))/2.057037k
 echo "Id"
 print -v(7)/2.078624k
 echo "Ic"
 print (v(5)-v(6))/3.092796k - (v(3)-v(2))/2.057037k
 
 print all
 .endc
 .end
