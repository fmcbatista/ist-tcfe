Circuito_t2

.INCLUDE ngspice_values.txt






.control
 op
 
 echo "Operating Point Analysis"
 
 print  V(6)-V(8) > Vx_p2.txt
 
 
 print all
 .endc
 .end
