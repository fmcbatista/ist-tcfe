Circuitot22

.INCLUDE ngspice2.txt

.INCLUDE Vxp2.tex

.control
 op
 
 echo "op2_TAB"
 print all
 print v(6)-v(8)
 print (v(6)-v(8))/vx#branch
 echo "op2_END"
 
 quit
 .endc
 .end
