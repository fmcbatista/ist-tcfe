Circuit_t2.3

.options savecurrents

.INCLUDE ngspice_3.txt


.ic v(6)=8.709810489  v(8)=0

.end

.control



op

echo "Transient Analysis"

tran 1e-6 20ms

plot v(6)

hardcopy trans.ps v(6)


.endc


.end
